
module canbacn_tb;
reg  [31:0]y,n;
wire [31:0]ketqua;
canbac_n u4(y,n,ketqua);
initial begin

y={32'b00111101010110000000000000000000}; //
n={32'b01000000100010000000000000000000}; // n
#100
y={32'b00111110010110000000000000000000}; 
n={32'b01000000010000000000000000000000}; //
#100
y={32'b01000000010110000000000000000000};	// 
n={32'b01000000100000000000000000000000}; //
#100
y={32'b00111111110110000000000000000000};	
n={32'b01000000010100000000000000000000}; // n =
#100
y={32'b01000000110010000000000000000000};
n={32'b01000000010000000000000000000000}; // n =
#100
y={32'b00111110010110000000000000000000};	
n={32'b01000000110000000000000000000000}; 
#100
y={32'b01000000110010000000000000000000};
n={32'b01000000011000100000000000000000}; // n =
#1000 $finish;
end 
endmodule
 
 