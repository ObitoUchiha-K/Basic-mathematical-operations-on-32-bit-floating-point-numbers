
module sinx_tb;
reg  [31:0]x;
wire [31:0]ketqua;
sin_x u4(x,ketqua);
initial begin
x={32'b11000000000000000000000000000000}; // -2
#300
x={32'b01000000010000000000000000000000}; // 3:
#300
x={32'b00111111010000000000000000000000}; // 0,75
#300
x={32'b00111111110110000000000000000000}; // 1,6875
#300
x={32'b00111111100000000000000000000000}; // 1
#300
x={32'b01000010111100000000000000000000}; // 120
#300
x={32'b11000011111001000000000000000000}; // -456
#300
x={32'b01000000110010010000111111011010}; // 2pi
#300
x={32'b00111111110010010000111111011010}; // pi/2
#300
x={32'b00000000000000000000000000000000}; // 0
#300
x={32'b00111100000000000000000000000000}; // 0,0078
#300
x={32'b00110001000000000000000000000000}; // ..10^-9
#300
x={32'b00110100000000000000000000000000}; //  ..10^-7
#300
x={32'b00111000000000000000000000000000}; // ..10^-5
#1000 $finish;
end 
endmodule


